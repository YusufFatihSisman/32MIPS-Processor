module and32(res, a, b);
	input [31:0] a, b;
	output [31:0] res;
	
	and a0(res[0], a[0], b[0]);
	and a1(res[1], a[1], b[1]);
	and a2(res[2], a[2], b[2]);
	and a3(res[3], a[3], b[3]);
	and a4(res[4], a[4], b[4]);
	and a5(res[5], a[5], b[5]);
	and a6(res[6], a[6], b[6]);
	and a7(res[7], a[7], b[7]);
	and a8(res[8], a[8], b[8]);
	and a9(res[9], a[9], b[9]);
	and a10(res[10], a[10], b[10]);
	and a11(res[11], a[11], b[11]);
	and a12(res[12], a[12], b[12]);
	and a13(res[13], a[13], b[13]);
	and a14(res[14], a[14], b[14]);
	and a15(res[15], a[15], b[15]);
	and a16(res[16], a[16], b[16]);
	and a17(res[17], a[17], b[17]);
	and a18(res[18], a[18], b[18]);
	and a19(res[19], a[19], b[19]);
	and a20(res[20], a[20], b[20]);
	and a21(res[21], a[21], b[21]);
	and a22(res[22], a[22], b[22]);
	and a23(res[23], a[23], b[23]);
	and a24(res[24], a[24], b[24]);
	and a25(res[25], a[25], b[25]);
	and a26(res[26], a[26], b[26]);
	and a27(res[27], a[27], b[27]);
	and a28(res[28], a[28], b[28]);
	and a29(res[29], a[29], b[29]);
	and a30(res[30], a[30], b[30]);
	and a31(res[31], a[31], b[31]);
	
endmodule