module alu32_testbench();
	reg [31:0] in1, in2;
	reg [2:0] aluCont;
	wire [31:0] result;
	wire [31:0] compareResult;
	wire zero;
	
	alu32 alu(result, compareResult, zero, in1, in2, aluCont);
	
	initial begin
	in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; aluCont = 3'b000;  
	#50;
	// and 00000000000000000000000000000111  11  
	in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; aluCont = 3'b001;  
	#50;
	// or 00100000000000000011000000011111   11
	in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; aluCont = 3'b010;  
	#50;
	// xor 00100000000000000011000000011000  11
	in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; aluCont = 3'b011;  
	#50;
	// add 00100000000000000011000000100110  11
	in1 = 32'b00000000000000000011000000011111; in2 = 32'b00100000000000000000000000000111; aluCont = 3'b111; 
	#50;
	// sub -011111111111111100111111101000  10

	in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; aluCont = 3'b000;
	#50;
	// and 00101000001001100001011001011110  11
	in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; aluCont = 3'b001;
	#50;
	// or 111110101111111101111111111111  11
	in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; aluCont = 3'b010;
	#50;
	// xor 110100101101100101101001101000  11
	in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; aluCont = 3'b011;
	#50;
	// add 100100011001001011001011001011101  11
	in1 = 32'b11111000011001110101111111011110; in2 = 32'b00101010101111100011011001111111; aluCont = 3'b111;
	#50;
	// sub 11001101101010010010100101011111  11


	in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; aluCont = 3'b000;
	#50;
	// and 00001111000011100011011000000000  11
	in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; aluCont = 3'b001;
	#50;
	// or 00111111111111110011111101111111  11
	in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; aluCont = 3'b010;
	#50;
	// xor 00110000111100010000100101111111  11
	in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; aluCont = 3'b011;
	#50;
	// add 1001111000011010111010101111111  11
	in1 = 32'b00001111000011110011111100011110; in2 = 32'b00111111111111100011011001100001; aluCont = 3'b111;
	#50;
	// sub -110000111011101111011101000011  10
	end
	 
	 
	initial begin
		$monitor("time = %2d, in1 = %32b, in2= %32b, alucont= %3b, result = %32b, compareResult = %32b, zero = %1b \n" , $time, in1, in2, aluCont, result, compareResult, zero);
	end
	 
 endmodule
